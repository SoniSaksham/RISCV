`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module memory(add,data_in,ALU_res,i_r,clk,rd_i,wr_rd,instr,data_out);
input [31:0]add,data_in,ALU_res;
input clk,rd_i,wr_rd,i_r;
output reg[31:0]instr;
output [31:0]data_out;
reg [31:0]rom[0:26];
reg [31:0]data[0:120];
wire [31:0]add1;

assign add1=i_r?ALU_res:add;

always@(posedge clk)
begin
if(rd_i)
instr<=rom[add];

if(wr_rd)
data[add1]<=data_in;
end
assign data_out=wr_rd?32'bz:data[add1];

initial
begin

rom[0]=32'h002082b3;
rom[1]=32'h402082b3;
rom[2]=32'h002092b3;
rom[3]=32'h0020a2b3;
rom[4]=32'h0020c2b3;
rom[5]=32'h0020d2b3;
rom[6]=32'h0020e2b3;
rom[7]=32'h4020d2b3;
rom[8]=32'h0020f2b3;
rom[9]=32'h00308293;
rom[10]=32'h0030a293;
rom[11]=32'h0030c293;
rom[12]=32'h0030e293;
rom[13]=32'h0030f293;
rom[14]=32'h0030a283;

rom[15]=32'h00309293; 

rom[16]=32'h0030d293;
rom[17]=32'h4030d293;
rom[18]=32'h0620a2a3;
rom[19]=32'h062082e3;
rom[20]=32'h062092e3;
rom[21]=32'h0620c2e3;
rom[22]=32'h0620d2e3;
rom[23]=32'h00c082e7;
rom[25]=32'h000082ef;
rom[26]=32'h000082b7;
rom[27]=32'h00008297;


data[0]=32'b00110010010101000011010000110111;
data[1]=32'b01110111010101000011010000010111;
data[2]=32'b11111111111111110101010001101111;
data[3]=32'b11110100010111110000010001100111;
data[4]=32'b10011010100011110000010001100011;
data[5]=32'b10111111011001000001010101100011;
data[6]=32'b10111100010101000100111001100011;
data[7]=32'b10111100010101000101011001100011;
data[8]=32'b10110010001100000110011001100011;
data[9]=32'b10011001001100000111011001100011;
data[10]=32'b11111011001100000000011000000011;
data[11]=32'b01100101001100000001011000000011;
data[12]=32'b11111010110111100010011000000011;
data[13]=32'b11111010110111100100011000000011;
data[14]=32'b11001010111011100101011000000011;
data[15]=32'b11001010111011100000011000100011;
data[16]=32'b11000111100011100001011000100011;
data[17]=32'b10011000011111100010011000100011;
data[18]=32'b10011000011111100000011000010011;
data[19]=32'b10010101011011100001011000010011;
data[20]=32'b11110100010011100010011000010011;
data[21]=32'b00110011010111100011011000010011;
data[22]=32'b00110011010100100100011000010011;
data[23]=32'b10010011010100100101011000010011;
data[24]=32'b11000000010100100110011000010011;
data[25]=32'b11001111010110000111011000010011;
data[26]=32'b00000000010110000001011000010011;
data[27]=32'b00000001010110000101011000010011;
data[28]=32'b01000001010110000101011000010011;
data[29]=32'b00000000010110000000011000110011;
data[30]=32'b01000000010110000000011000110011;
data[31]=32'b00000000010110000001011000110011;
data[32]=32'b00000000111110000010011000110011;
data[33]=32'b00000000111111110011011000110011;
data[34]=32'b00000000100110010100011000110011;
data[35]=32'b00000000111110010101011000110011;
data[36]=32'b01000000111110010101011000110011;
data[37]=32'b00000000111110010110011000110011;
data[38]=32'b00000000111110010111011000110011;
data[39]=32'b10011000011111100000011000010011;
data[108]=32'b10011000011111100000011000010011;

end
endmodule




